// =============================================================
// sigmoid_lut.v — Sigmoid Activation LUT
// =============================================================
// 256-entry lookup table implementing sigmoid(x) = 1/(1+e^-x)
//
// Input  : 8-bit index (taken from bits [14:7] of Q4.12 accumulator)
// Output : Q4.12 sigmoid value (range 0.0 to 1.0)
//
// Index mapping:
//   index 0   → input = -8.0  → sigmoid ≈ 0.000335
//   index 128 → input =  0.0  → sigmoid = 0.5
//   index 255 → input = +7.9375 → sigmoid ≈ 0.99966
//
// To use: addr = accumulator[14:7]
//   (takes integer part + top 3 fractional bits of Q4.12 value)
// =============================================================

module sigmoid_lut (
    input  wire        clk,
    input  wire [7:0]  addr,   // 8-bit index
    output reg  [15:0] data    // Q4.12 sigmoid output
);
    // 256 x 16-bit ROM — synthesizes to LUTRAM or BRAM on Xilinx
    reg [15:0] lut [0:255];

    // Load precomputed Q4.12 values generated by weight_extractor.py
    initial $readmemh("sigmoid_lut.hex", lut);

    // Registered output — 1 clock cycle latency
    always @(posedge clk)
        data <= lut[addr];

endmodule
